`timescale 1ns/100ps
module rem_tb ();
reg [2:0] A;
reg [2:0] B;
wire [2:0] R;
wire DZF;
wire ZF;
wire SF;
integer f;
rem test (.A(A),
.B(B),
.R(R),
.DZF(DZF),
.SF(SF),
.ZF(ZF));
initial begin
    f = $fopen("rem.txt","w");
    A[1:0]=2'b00; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b0; #10;    
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b0; #10;   
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b1; #10;    
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b10; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b01; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b00; A[2]=1'b0; B[2]=1'b1; #10;   
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b11; A[2]=1'b0; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b0; #10;    
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b0; #10;   
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b0; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b00; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b1; #10;    
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b01; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b10; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b10; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b01; A[2]=1'b1; B[2]=1'b1; #10;
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b00; A[2]=1'b1; B[2]=1'b1; #10;   
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    A[1:0]=2'b11; B[1:0]=2'b11; A[2]=1'b1; B[2]=1'b1; #10;    
    $fdisplay(f,"A = %03b ,B= %03b ,R = %03b,DZF = %0b,SF = %0b,ZF = %0b",A,B,R,DZF,SF,ZF);
    $fclose(f);
end
endmodule